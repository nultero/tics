module tics

